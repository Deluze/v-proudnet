module proud

// todo: can't use enum as generic even if marked as u8..
struct HostIDArray {
	CFastArray[u8]
}