module proud

struct HostIDArray {
	CFastArray[HostID]
}