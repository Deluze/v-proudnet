module proud

struct HostIDArray {

}
