module main

import net
import proud

fn main() {
}
