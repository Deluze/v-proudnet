module proud

type HostIDArray = CFastArray[HostID]