module proud

struct CNetServer {
	CoreEventFunctions
}